-- Test Bench for Counter.
library IEEE;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;



entity tb_bs is
  GENERIC (n : INTEGER :=4 ;m : INTEGER :=3);
end tb_bs;

architecture rtl of tb_bs is  
COMPONENT BarrelShfter IS
  GENERIC (n : INTEGER;m : INTEGER);
  PORT (    x: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
			yi: IN STD_LOGIC_VECTOR (n-1 DOWNTO 0);
            s: OUT STD_LOGIC_VECTOR(n-1 downto 0));
END COMPONENT;

signal  x:STD_LOGIC_VECTOR (n-1 DOWNTO 0);
signal	yi :STD_LOGIC_VECTOR (n-1 DOWNTO 0);
signal	s :STD_LOGIC_VECTOR(n-1 downto 0);

begin
        tester : BarrelShfter generic map (n=>n,m=>m) port map(
			x=>x,yi=>yi,s=>s
		);
        
        testbench : process
        begin
          --------- start of stimulus section - ver1 ------------------
          x <="1111";
		   yi <="0000";
		   for i in 0 to 4 loop
			wait for 50 ns;
			yi <= yi +1;
		  end loop;
          --------- end of stimulus section----------------------------
		  wait;
        end process testbench;
        
end rtl;
